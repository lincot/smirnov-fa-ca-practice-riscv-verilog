module xor4(input logic x0, x1, x2, x3, output logic y);
    assign y = x0 ^ x1 ^ x2 ^ x3;
endmodule